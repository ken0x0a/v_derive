module common

import v.ast { EnumDecl, Stmt, StructDecl, SumTypeDecl }
import v.token
import codegen { Codegen }
import util { get_type_name_without_module }

// ```v
// pub fn (self ItemB) bin_len() int {
// 	mut len := 0
// 	len += bincode.len(self.b)
// 	len += bincode.len(self.bb)
// 	len += bincode.len(self.bbb)
// 	return len
// }
// ```
pub fn add_len_fn_for_struct(mut cg Codegen, decl StructDecl) {
	fn_name := common.fn_method_name_len
	mut params := []ast.Param{cap: decl.fields.len}
	// return_type := cg.find_type_or_add_placeholder(get_type_name_without_module(decl.name),
	// 	.v)

	mut body_stmts := []Stmt{cap: decl.fields.len + 2}
	body_stmts << base_assign_stmt(mut cg)
	for field in decl.fields {
		body_stmts << gen_plus_assign_len_call(mut cg, field)
	}
	body_stmts << Stmt(ast.Return{
		exprs: [cg.ident(common.ident_name_len)]
	})
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: ast.int_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}

// ```v
// len += bincode.len(self.b)
// ```
fn gen_plus_assign_len_call(mut cg Codegen, field ast.StructField) ast.Stmt {
	field_name := field.name

	field_sel := ast.SelectorExpr{ // 'self.$field'
		field_name: field_name
		expr: cg.ident(ident_name_self)
		scope: cg.scope()
	}

// TODO: handle type here `array` `map` & ...
	right := get_call_len(mut cg, field, field_sel)

	return ast.AssignStmt{
		left: [cg.ident(ident_name_len)]
		right: [right]
		op: token.Kind.plus_assign
	}
}

// ```v
// bincode.len(self.b)
// ```
fn get_call_len(mut cg Codegen, field ast.StructField, sel ast.Expr) ast.Expr {
	return ast.CallExpr{
		name: 'len'
		left: cg.ident(mod_name)
		args: [
			ast.CallArg{
				expr: sel
			}
		]
		scope: cg.scope()
		is_method: true
	}
}