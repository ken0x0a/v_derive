module common

import v.ast { EnumDecl, Stmt, StructDecl, SumTypeDecl }
import v.token
import term
import codegen { Codegen }
import util { get_type_name_without_module }

const (
	macro_name                 = 'BinEncode'
	mod_name                   = 'bincode'
	const_str_0_bytes_for_len  = 'num_bytes_for_len'
	bytes_len_int              = 4
	fn_method_name_len         = 'bin_len'
	fn_method_name_encode      = 'bin_encode'
	fn_method_name_encode_self = 'bin_encode_self'
	fn_method_name_decode      = 'bin_decode'
	ident_name_len             = 'len'
	ident_name_self            = 'self'
)

pub fn get_fn_name_decode(name string) string {
	base := util.to_snake_case(get_type_name_without_module(name))
	return 'bin_decode__$base'
}

fn base_assign_stmt(mut cg Codegen) Stmt {
	return Stmt(ast.AssignStmt{
		left: [cg.ident_opt(common.ident_name_len, is_mut: true)]
		right: [cg.integer_literal(0)]
		op: token.Kind.decl_assign
	})
}


// ```v
// pub fn (self OneOf) bin_len() int {
// 	mut len := 0
// 	len += bincode.len_for<byte>()
// 	len += match self {
// 		ItemA { self.bin_len() }
// 		ItemB { self.bin_len() }
// 	}
// 	return len
// }
// ```
pub fn add_len_fn_for_sumtype(mut cg Codegen, decl SumTypeDecl) {
	fn_name := common.fn_method_name_len
	mut params := []ast.Param{}

	mut body_stmts := []Stmt{cap: decl.variants.len + 5}
	body_stmts << base_assign_stmt(mut cg)
	body_stmts << plus_assign_sumtype_type(mut cg)
	body_stmts << plus_assign_sumtype_match(mut cg, decl)
	body_stmts << Stmt(ast.Return{
		exprs: [cg.ident(common.ident_name_len)]
	})

	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: ast.int_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}

// ```v
// pub fn (self ItemB) bin_len() int {
// 	mut len := 0
// 	len += bincode.len(self.b)
// 	len += bincode.len(self.bb)
// 	len += bincode.len(self.bbb)
// 	return len
// }
// ```
pub fn add_len_fn_for_struct(mut cg Codegen, decl StructDecl) {
	fn_name := common.fn_method_name_len
	mut params := []ast.Param{cap: decl.fields.len}
	// return_type := cg.find_type_or_add_placeholder(get_type_name_without_module(decl.name),
	// 	.v)

	mut body_stmts := []Stmt{cap: decl.fields.len + 2}
	body_stmts << base_assign_stmt(mut cg)
	for field in decl.fields {
		body_stmts << set_value_stmt_or_skip(mut cg, field)
	}
	body_stmts << Stmt(ast.Return{
		exprs: [cg.ident(common.ident_name_len)]
	})
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: ast.int_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}

// Enum value is always `int` => 4 bytes in Vlang
// Generates:
//
// ```v
// [inline]
// fn (self EnumName) bin_len() int {
// 	return 4
// }
// ```
pub fn add_len_fn_for_enum(mut cg Codegen, decl EnumDecl) {
	fn_name := common.fn_method_name_len
	params := []ast.Param{}
	return_type := ast.int_type
	mut body_stmts := []Stmt{}

	body_stmts << Stmt(ast.Return{
		exprs: [
			cg.integer_literal(common.bytes_len_int),
		]
	})
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: return_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}
