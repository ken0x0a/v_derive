module deser_json

import v.ast
import v.token
import tool.codegen.codegen { Codegen }

fn get_map_depth(type_name string) int {
	mut temp := type_name
	mut depth := 0
	for {
		if temp.starts_with('map[string]') {
			depth += 1
			temp = temp[10..]
		} else {
			return depth
		}
	}
	return depth
}

fn register_map_fn_if_not_exist(mut self Codegen, typ ast.Type, typ_arg string, fn_name string, depth int) {
	if fn_name in self.table.fns {
		eprintln('"$fn_name" is already registered')
	} else {
		typ_sym := self.table.sym(typ)
		body_stmts := [
			// obj := j.as_map()
			ast.Stmt(ast.AssignStmt{
				left: [self.ident(json2_map_name)]
				right: [ast.Expr(ast.CallExpr{
					name: 'as_map'
					left: self.ident(json2_any_param_name)
					scope: self.scope()
					is_method: true
				})]
				op: token.Kind.decl_assign // op: token.Kind.and // op: token.Kind.assign
			}),
			// 
			ast.Stmt(ast.AssignStmt{
				left: [self.ident_opt('res', is_mut: true)]
				right: [ast.Expr(ast.MapInit{
					typ: typ
				})]
				op: token.Kind.decl_assign // op: token.Kind.and // op: token.Kind.assign
			}),
			// ast.Stmt(ast.AssignStmt{
			// 	left: [self.ident(json2_map_name)]
			// 	right: [
			// 		ast.Expr(ast.CallExpr{
			// 			name: 'as_map'
			// 			left: self.ident('j')
			// 			scope: self.scope()
			// 			is_method: true
			// 		})
			// 	]
			// 	// op: token.Kind.assign
			// 	op: token.Kind.decl_assign
			// 	// op: token.Kind.and
			// })
			ast.ForInStmt{
				key_var: 'key'
				val_var: 'val'
				cond: self.ident(json2_map_name)
				scope: self.scope()
				stmts: [
					ast.Stmt(ast.AssignStmt{
					left: [
						ast.Expr(ast.IndexExpr{
							index: self.ident('key')
							left: self.ident('res')
						}),
					]
					right: [
						ast.Expr(ast.CallExpr{
							name: if depth == 1 {
								get_decode_fn_name(typ_arg)
							} else {
								get_decode_map_fn_name(typ_arg, depth - 1)
							}
							args: [ast.CallArg{
								expr: self.ident('val')
							}]
							scope: self.scope()
							is_method: false
							or_block: ast.OrExpr{
								kind: .propagate
							}
						}),
					]
					// op: token.Kind.assign
					op: token.Kind.assign
					// op: token.Kind.and
				}),
				]
			},
			ast.Return{
				exprs: [self.ident('res')]
			},
		]

		// return_type := self.find_type_or_add_placeholder(typ_sym.name, .v)
		return_type := typ.set_flag(.optional)
		$if debug_ast ? {
			dump(self.find_type_or_add_placeholder('map[string]json2.Any', .v))
			dump(typ)
		}
		params := [ast.Param{
			name: json2_any_param_name
			typ: self.find_type_or_add_placeholder('json2.Any', .v)
		}]

		// ## Register to table
		fn_def := ast.Fn{
			name: fn_name
			params: params
			return_type: return_type
		}
		// self.table.fns[fn_name] = fn_def

		self.add_fn(
			name: fn_name
			return_type: return_type
			body_stmts: body_stmts
			params: params
			comments: [self.gen_comment(text: 'generated by macro "derive_Deser')]
		)
		self.table.find_or_register_fn_type(typ_sym.mod, fn_def, false, true)
	}
}
