module de

import v.ast {Stmt}
import v.token
import codegen { Codegen }
import common
import util {get_type_name_without_module}

pub const (
	macro_name = 'DeserBin'
)
const (
	ident_name_bytes = 'b'
	ident_name_decoded_len = 'd_len'
	ident_name_decode_pos = 'pos'
)

// ```v
// mut pos := 0
// ```
fn base_assign_stmt(mut cg Codegen) Stmt {
	return Stmt(ast.AssignStmt{
		left: [cg.ident_opt(ident_name_decode_pos, is_mut: true)]
		right: [cg.integer_literal(0)]
		op: token.Kind.decl_assign
	})
}
// ```v
// defer {
// 	d_len += pos
// }
// ```
fn gen_defer_stmt(mut cg Codegen) ast.DeferStmt {
	return ast.DeferStmt{
		stmts: [ast.Stmt(ast.AssignStmt{
			left: [cg.ident(ident_name_decoded_len)]
			right: [cg.ident(ident_name_decode_pos)]
			op: token.Kind.plus_assign
		})]
	}
}

// ```v
// name: bincode.decode<string>(buf, mut pos)
// ```
fn gen_struct_init_field(mut cg Codegen, field ast.StructField, idx int) ast.StructInitField {
	arg1 := if idx == 0 {
		ast.CallArg{
			expr: cg.ident(ident_name_bytes)
		}
	} else {
		ast.CallArg{
			expr: ast.IndexExpr{
				left: cg.ident(ident_name_bytes)
				index: ast.RangeExpr{has_low: true, low: cg.ident(ident_name_decode_pos)}
			}
		}
	}
	return ast.StructInitField{
		name: field.name
		expr: ast.CallExpr{
			name: 'decode',
			left: cg.ident(common.mod_name)
			scope: cg.scope()
			is_method: true
			concrete_types: [field.typ]
			args: [arg1, ast.CallArg{
				expr: cg.ident(ident_name_decode_pos)
				is_mut: true
			}]
		}
	}
}
// generates
// ```vlang
// fn bin_decode__product(buf []byte, mut d_len &int) Product {
// 	mut pos := 0
// 	defer {
// 		d_len += pos
// 	}
// 	return Product{
// 		name: bincode.decode<string>(buf, mut pos)
// 		desc: bincode.decode<string>(buf[pos..], mut pos)
// 		inventory: bincode.decode<u32>(buf[pos..], mut pos)
// 		price: bincode.decode<f64>(buf[pos..], mut pos)
// 	}
// }
// ```
pub fn add_decode_fn_for_struct(mut cg Codegen, decl ast.StructDecl) {
	fn_name := common.get_fn_name_decode(decl.name)
	mut params := get_params(mut cg)
	return_type := cg.find_type_or_add_placeholder(get_type_name_without_module(decl.name), .v)
	typ_sym := cg.table.find_sym(decl.name) or {panic(err)}

	mut body_stmts := []Stmt{cap: decl.fields.len + 3}
	body_stmts << base_assign_stmt(mut cg)
	defer_stmt := gen_defer_stmt(mut cg)
	body_stmts << defer_stmt
	mut fields := []ast.StructInitField{ cap: decl.fields.len}
	for idx, field in decl.fields {
		fields << gen_struct_init_field(mut cg, field, idx)
	}
	body_stmts << Stmt(ast.Return{
		exprs: [ast.Expr(ast.StructInit{
			typ: return_type
			fields: fields
		})]
	})
	// ## Register to table
	fn_def := ast.Fn{
		name: fn_name
		params: params
		return_type: return_type
	}

	cg.add_fn(
		name: fn_name
		return_type: return_type
		body_stmts: body_stmts
		params: params
		is_pub: true
		comments: [cg.gen_comment(text: 'generated by macro "$macro_name"')]
	)
	cg.table.find_or_register_fn_type(typ_sym.mod, fn_def, false, true)
}
pub fn add_decode_method_for_struct(mut cg Codegen, decl ast.StructDecl) {
	fn_name := common.get_fn_name_decode(decl.name)
	mut params := []ast.Param{cap: decl.fields.len}
	// return_type := cg.find_type_or_add_placeholder(get_type_name_without_module(decl.name), .v)

	mut body_stmts := []Stmt{cap: decl.fields.len + 2}
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: ast.int_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}
