module common

import v.ast {Stmt, EnumDecl}
import codegen { Codegen }

// Enum value is always `int` => 4 bytes in Vlang
// Generates:
//
// ```v
// [inline]
// fn (self EnumName) bin_len() int {
// 	return 4
// }
// ```
pub fn add_len_fn_for_enum(mut cg Codegen, decl EnumDecl) {
	fn_name := common.fn_method_name_len
	params := []ast.Param{}
	return_type := ast.int_type
	mut body_stmts := []Stmt{}

	body_stmts << Stmt(ast.Return{
		exprs: [
			cg.integer_literal(common.bytes_len_int),
		]
	})
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: return_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$common.macro_name"'),
		]
	)
}
