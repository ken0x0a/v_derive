module as_map

import v.ast
import v.token
import term
import tool.codegen.codegen { Codegen }

pub const (
	name_as_http_params    = 'AsHttpParams'
	fn_name_as_http_params = 'as_http_params'
)
const (
	json2_map_name         = 'obj'
)

// generates
// ```vlang
// fn (mut self Struct) as_http_params() map[string]string {
// 	mut obj := map[string]string{}
// 	obj['name'] = self.name
// 	obj['f64_val'] = f64(self.f64_val).str().trim_right('.') // as str
// 	return obj
// }
// ```
pub fn add_as_http_params_fn_for_struct(mut self Codegen, stmt ast.StructDecl) {
	mut body_stmts := []ast.Stmt{}
	return_type := self.find_type_or_add_placeholder('map[string]string', .v)
	body_stmts << ast.Stmt(ast.AssignStmt{
		left: [self.ident_opt(json2_map_name, is_mut: true)]
		right: [
			ast.Expr(ast.MapInit{
				typ: return_type
			})
		]
		op: token.Kind.decl_assign
	})

	for field in stmt.fields {
		js_field_name := get_js_field_name(field)
		body_stmts << set_value_stmt(mut self, field.name, js_field_name, field.typ)
	}

	body_stmts << ast.Stmt(ast.Return{
		exprs: [self.ident(json2_map_name)]
	})
	self.add_struct_method(
		struct_name: stmt.name.split('.').last()
		is_mut: false
		name: fn_name_as_http_params
		return_type: return_type
		body_stmts: body_stmts
		params: []
		comments: [
			self.gen_comment(text: 'generated by derive macro "AsHttpParams'),
			self.gen_comment(text: 'Example: $fn_name_as_http_params'),
		]
	)
}

fn set_value_stmt(mut self Codegen, field_name string, js_field_name string, typ ast.Type) ast.Stmt {
	field := ast.SelectorExpr{ // 'self.field'
		field_name: field_name
		expr: self.ident('self')
		scope: self.scope()
	}
	right := if typ == ast.string_type {
		ast.Expr(field)
	} else if self.table.get_type_symbol(typ).has_method('str') {
		mut type_sym := self.table.get_type_symbol(typ)
		print(field_name)
		dump(type_sym.name)

		ast.Expr(ast.CallExpr{
			name: 'str'
			left: field
			scope: self.scope()
			is_method: true
		})
	} else {
		mut type_sym := self.table.get_type_symbol(typ)
		info := type_sym.info
		// ISSUE: https://github.com/vlang/v/issues/9419
		_ := match info {
			ast.Alias {
				type_sym = self.table.get_type_symbol(info.parent_type)
				_ = $if debug {
					println(term.red(type_sym.name))
					dump(type_sym.name)
					true
				} $else {
					true
				}
				true // ISSUE: 9419
			}
			else {true} // ISSUE: 9419
		}
		// if info is ast.Alias {
		// 	type_sym = self.table.get_type_symbol(info.parent_type)
		// 	println(term.red(type_sym.name))
		// 	dump(type_sym.name)
		// }

		// dump(field_name)
		// dump(type_sym.name)
		// dump(type_sym.methods)
		// dump(type_sym.info)
		match type_sym.info {
			ast.Map {
				ast.Expr(field)
			}
			ast.Array {
				// field.map(it.str()).join('')
				ast.Expr(ast.CallExpr{
					name: 'join'
					args: [ast.CallArg{ expr: self.string_literal('') }]
					left: ast.CallExpr{
						name: 'map'
						args: [ast.CallArg {
							expr: ast.CallExpr{
								name: 'str'
								left: self.ident('it')
								scope: self.scope()
								is_method: true
							}
						}]
						left: field
						scope: self.scope()
						is_method: true
					}
					scope: self.scope()
					is_method: true
				})
			}
			ast.Enum {
				ast.Expr(ast.CallExpr{
					name: 'str'
					left: field
					scope: self.scope()
					is_method: true
				})
			}
			else {
				// print('${field_name:-20}')
				// dump(type_sym.name)

				ast.Expr(ast.CallExpr{
					name: 'str'
					left: field
					scope: self.scope()
					is_method: true
				})
			}
		}
	}
	return ast.AssignStmt{
		left: [ast.Expr(ast.IndexExpr{
			index: self.string_literal(js_field_name)
			left: self.ident(json2_map_name)
		})]
		right: [right]
		op: token.Kind.assign
	}
}

fn get_js_field_name(field ast.StructField) string {
	mut name := field.name
	for attr in field.attrs {
		if attr.name == 'json' {
			name = attr.arg
		}
		$if debug_attr ? {
			println(attr)
		}
	}
	return name
}
