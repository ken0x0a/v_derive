module de

import v.ast { Stmt }
import v.token
import codegen { Codegen }
import common
import util { get_type_name_without_module }

// generates
// ```vlang
// fn bin_decode__one_of(buf []u8, mut d_len &int) OneOf {
// 	mut pos := 0
// 	typ := decode<u8>(buf, mut pos)
// 	defer {
// 		d_len += pos
// 	}
// 	match typ {
// 		1 { return OneOf(bin_decode__item_a(buf[pos..], mut pos)) }
// 		2 { return OneOf(bin_decode__item_b(buf[pos..], mut pos)) }
// 		else { panic('Unsupported type `$typ`') }
// 	}
// }
// ```
pub fn add_decode_fn_for_sumtype_fn(mut cg Codegen, decl ast.SumTypeDecl) {
	fn_name := common.get_fn_name_decode(decl.name)
	mut params := get_params(mut cg)
	return_type := cg.find_type_or_add_placeholder(get_type_name_without_module(decl.name),
		.v)
	typ_sym := cg.table.find_sym(decl.name) or { panic(err) }

	mut body_stmts := []Stmt{cap: decl.variants.len + 2}
	body_stmts << base_assign_stmt(mut cg)
	defer_stmt := gen_defer_stmt(mut cg)
	body_stmts << defer_stmt
	ident_typ := cg.ident('typ')
	body_stmts << ast.AssignStmt{
		left: [ident_typ]
		right: [
			ast.Expr(ast.CallExpr{
				name: 'decode'
				left: cg.ident(common.mod_name)
				scope: cg.scope()
				is_method: true
				concrete_types: [ast.u8_type]
				args: [ast.CallArg{
					expr: cg.ident(ident_name_bytes)
				}, ast.CallArg{
					expr: cg.ident(ident_name_decode_pos)
					is_mut: true
				}]
			}),
		]
		op: token.Kind.decl_assign
	}
	body_stmts << ast.ExprStmt{
		expr: gen_sumtype_match_expr(mut cg, decl, return_type)
	}

	// ## Register to table
	fn_def := ast.Fn{
		name: fn_name
		params: params
		return_type: return_type
	}

	cg.add_fn(
		name: fn_name
		return_type: return_type
		body_stmts: body_stmts
		params: params
		is_pub: true
		comments: [cg.gen_comment(text: 'generated by macro "$macro_name"')]
	)
	cg.table.find_or_register_fn_type(typ_sym.mod, fn_def, false, true)
}

// ```v
// match typ {
// 	1 { return OneOf(bin_decode__item_a(buf[pos..], mut pos)) }
// 	2 { return OneOf(bin_decode__item_b(buf[pos..], mut pos)) }
// 	else { panic('Unsupported type `$typ`') }
// }
// ```
fn gen_sumtype_match_expr(mut cg Codegen, decl ast.SumTypeDecl, return_type ast.Type) ast.Expr {
	mut branches := []ast.MatchBranch{cap: decl.variants.len}
	for idx, var in decl.variants {
		sym := cg.table.sym(var.typ)
		fn_name := common.get_fn_name_decode(sym.name)

		branches << ast.MatchBranch{
			scope: cg.scope()
			exprs: [cg.integer_literal(idx + 1)]
			stmts: [
				Stmt(ast.Return{
					exprs: [
						ast.Expr(ast.CastExpr{
							typ: return_type
							expr: ast.CallExpr{
								name: fn_name
								scope: cg.scope()
								args: [
									ast.CallArg{
										expr: ast.IndexExpr{
											left: cg.ident(ident_name_bytes)
											index: ast.RangeExpr{
												has_low: true
												low: cg.ident(ident_name_decode_pos)
											}
										}
									},
									ast.CallArg{
										expr: cg.ident(ident_name_decode_pos)
										is_mut: true
									},
								]
							}
						}),
					]
				}),
			]
		}
	}
	branches << ast.MatchBranch{
		scope: cg.scope()
		is_else: true
		stmts: [
			Stmt(ast.ExprStmt{
				expr: ast.CallExpr{
					name: 'panic'
					scope: cg.scope()
					args: [
						ast.CallArg{
							expr: cg.string_literal('Unsupported type `\$typ` < $decl.variants.len')
						},
					]
				}
			}),
		]
	}
	return ast.Expr(ast.MatchExpr{
		is_expr: true
		return_type: return_type
		cond: cg.ident('typ')
		branches: branches
	})
}
