module ser

import v.ast
import v.pref
import v.parser
import codegen

fn test_enum_bin_encode() ? {
	test_text := '
enum TestEnum {
	a
	b
	c
}
'
	mut table := ast.new_table()
	// parsed := parser.parse_file(filename, table, .parse_comments, &pref.Preferences{})
	// mut gen := codegen.new_with_table(mod_name: module_name, table: table)
	mut gen := codegen.new_with_table(table: table)
	parsed := parser.parse_text(test_text, 'dummy.v', gen.table, .parse_comments, &pref.Preferences{})
	module_name := parsed.mod.name.split('.').last()
	println('module_name: $module_name ($parsed.mod.name)')
	dump(parsed.stmts)
	assert parsed.stmts.len == 2
	assert parsed.stmts[1] is ast.EnumDecl
	add_encode_fn_for_enum(mut gen, parsed.stmts[1] as ast.EnumDecl)
	dump(gen)
	assert gen.to_code_string() == 'module main

// generated by macro "BinEncode"
pub fn (self TestEnum) bin_encode(mut b []u8) int {
	return unsafe { bincode.encode(int(self)) }
}
'
}

fn test_struct_bin_encode() ? {
	test_text := '
struct Test {
	a int
	b string
	c u64
}
'
	mut table := ast.new_table()
	// parsed := parser.parse_file(filename, table, .parse_comments, &pref.Preferences{})
	// mut gen := codegen.new_with_table(mod_name: module_name, table: table)
	mut gen := codegen.new_with_table(table: table)
	parsed := parser.parse_text(test_text, 'dummy.v', gen.table, .parse_comments, &pref.Preferences{})
	module_name := parsed.mod.name.split('.').last()
	println('module_name: $module_name ($parsed.mod.name)')
	dump(parsed.stmts)
	assert parsed.stmts.len == 2
	assert parsed.stmts[1] is ast.StructDecl
	add_encode_fn_for_struct(mut gen, parsed.stmts[1] as ast.StructDecl)
	// dump(gen)
	expected := 'module main

// generated by macro "SerBin"
pub fn (self Test) bin_encode(mut b []u8) int {
	mut pos := 0
	pos += bincode.encode(mut b, self.a)
	pos += bincode.encode(mut b[pos..], self.b)
	pos += bincode.encode(mut b[pos..], self.c)
	return pos
}
'
	result := gen.to_code_string()
	// for i in 0..expected.len {
	// 	println(i)

	// 	assert result[i] == expected[i]
	// }
	// assert result.len == expected.len
	assert result == expected
}

fn test_sumtype_bin_encode() ? {
	test_text := '
type OneOf = ItemA | ItemB
struct ItemA {
	a int
}
struct ItemB {
	b string
}
'
	mut table := ast.new_table()
	// parsed := parser.parse_file(filename, table, .parse_comments, &pref.Preferences{})
	// mut gen := codegen.new_with_table(mod_name: module_name, table: table)
	mut gen := codegen.new_with_table(table: table)
	parsed := parser.parse_text(test_text, 'dummy.v', gen.table, .parse_comments, &pref.Preferences{})
	module_name := parsed.mod.name.split('.').last()
	println('module_name: $module_name ($parsed.mod.name)')
	assert parsed.stmts.len == 4
	assert parsed.stmts[1] is ast.TypeDecl
	add_encode_fn_for_sumtype(mut gen, parsed.stmts[1] as ast.TypeDecl as ast.SumTypeDecl)
	dump(gen.file.stmts)
	assert gen.to_code_string() == 'module main

// generated by macro "SerBin"
pub fn (self OneOf) bin_encode(mut b []u8) int {
	mut pos := 0
	pos += match self {
		ItemA {
			pos += unsafe { bincode.encode<u8>(mut b, 1) }
			unsafe { bincode.encode(mut b[pos..], self) }
		}
		ItemB {
			pos += unsafe { bincode.encode<u8>(mut b, 2) }
			unsafe { bincode.encode(mut b[pos..], self) }
		}
	}
	return pos
}
'
}
