module common

import v.ast { Stmt, SumTypeDecl }
import v.token
import codegen { Codegen }
import util

// ```v
// pub fn (self OneOf) bin_len() int {
// 	mut len := 0
// 	len += bincode.len_for<u8>()
// 	len += match self {
// 		ItemA { self.bin_len() }
// 		ItemB { self.bin_len() }
// 	}
// 	return len
// }
// ```
pub fn add_len_fn_for_sumtype(mut cg Codegen, decl SumTypeDecl) {
	fn_name := fn_method_name_len
	mut params := []ast.Param{}

	mut body_stmts := []Stmt{cap: decl.variants.len + 5}
	body_stmts << base_assign_stmt(mut cg)
	body_stmts << plus_assign_sumtype_type(mut cg)
	body_stmts << plus_assign_sumtype_match(mut cg, decl)
	body_stmts << Stmt(ast.Return{
		exprs: [cg.ident(ident_name_len)]
	})

	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: ast.int_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$macro_name"'),
		]
	)
}

// ```v
// len += bincode.len_for<u8>()
// ```
fn plus_assign_sumtype_type(mut cg Codegen) Stmt {
	right := ast.Expr(ast.CallExpr{
		name: 'len_for'
		concrete_types: [ast.byte_type]
		left: cg.ident(mod_name)
		scope: cg.scope()
		is_method: true
	})
	return ast.AssignStmt{
		left: [cg.ident(ident_name_len)]
		right: [right]
		op: token.Kind.plus_assign
	}
}

// ```v
// len += match self {
// 	ItemA { self.bin_len() }
// 	ItemB { self.bin_len() }
// }
// ```
fn plus_assign_sumtype_match(mut cg Codegen, decl SumTypeDecl) Stmt {
	mut branches := []ast.MatchBranch{cap: decl.variants.len}
	for var in decl.variants {
		sym := cg.table.sym(var.typ)
		dump(sym.info)
		branches << ast.MatchBranch{
			scope: cg.scope()
			exprs: [cg.ident(util.get_type_name_without_module(sym.name))]
			stmts: [
				Stmt(ast.ExprStmt{
					expr: ast.CallExpr{
						name: fn_method_name_len
						left: cg.ident(ident_name_self)
						scope: cg.scope()
						is_method: true
					}
				}),
			]
		}
	}
	right := ast.Expr(ast.MatchExpr{
		is_expr: true
		return_type: ast.string_type
		cond: cg.ident('self')
		branches: branches
	})
	return ast.AssignStmt{
		left: [cg.ident(ident_name_len)]
		right: [right]
		op: token.Kind.plus_assign
	}
}
