module ser_json

import v.ast
import v.token
import term
import tool.codegen.codegen { Codegen }

pub const (
	macro_name = 'Ser_json'
)
const (
	json2_map_name            = 'obj'
	json2_any_param_name      = 'j'
	encode_json_pub_fn_prefix = 'ser_json'
	encode_json_member_name   = 'to_json'
	encode_json_fn_name       = 'macro_ser_json'
	encode_json_fn_arg_name   = 'src'
	encode_json_map_fn_name   = 'macro_ser_json_map'
	encode_json_array_fn_name = 'macro_ser_json_array'
)

// generates
// ```vlang
// fn (self Struct) to_json() string {
// 	mut obj := map[string]json2.Any{}
// 	obj['name'] = self.name
// 	obj['f64_val'] = f64(self.f64_val).str().trim_right('.') // as str
// 	return obj.str()
// }
// ```
pub fn add_encode_json(mut self Codegen, stmt ast.StructDecl) {
	// mut body_stmts := []ast.Stmt{}
	mut body_stmts := get_encode_json_base_stmts(mut self)
	for field in stmt.fields {
		js_field_name := get_js_field_name(field)
		body_stmts << set_value_stmt(mut self, field.name, js_field_name, field.typ)
	}
	body_stmts << ast.Stmt(
		ast.Return{
			exprs: [ast.Expr(
				ast.CallExpr{
					name: 'str'
					left: self.ident(json2_map_name)
					scope: self.scope()
					is_method: true
				}
			)]
		}
	)
	self.add_struct_method(
		struct_name: stmt.name.split('.').last()
		is_mut: false
		name: ser_json.encode_json_member_name
		return_type: ast.string_type
		body_stmts: body_stmts
		params: []
		comments: [
			self.gen_comment(text: 'generated by macro "derive_Deser'),
			self.gen_comment(
				text: 'Example: $ser_json.encode_json_fn_name<${stmt.name.split('.').last()}>(text)'
			),
		]
	)
}

// mut obj := map[string]json2.Any{}
fn get_encode_json_base_stmts(mut self Codegen) []ast.Stmt {
	return [
		ast.Stmt(ast.AssignStmt{
			left: [self.ident_opt(ser_json.json2_map_name, is_mut: true)]
			right: [
				ast.Expr(ast.MapInit{
					typ: self.find_type_or_add_placeholder('map[string]json2.Any', .v)
				})
			]
			op: token.Kind.decl_assign
		}),
	]
}

fn set_value_stmt(mut self Codegen, field_name string, js_field_name string, typ ast.Type) ast.Stmt {
	field := ast.SelectorExpr{ // 'self.field'
		field_name: field_name
		expr: self.ident('self')
		scope: self.scope()
	}

	right := get_type_recursively(mut self, field, typ)

	return ast.AssignStmt{
		left: [ast.Expr(ast.IndexExpr{
			index: self.string_literal(js_field_name)
			left: self.ident(ser_json.json2_map_name)
		})]
		right: [right]
		op: token.Kind.assign
	}
}
fn get_type_recursively(mut self Codegen, field ast.Expr, typ ast.Type) ast.Expr {
	// fallback to parent type, if type has no `str` method
	mut type_sym := self.table.get_type_symbol(typ)
	if type_sym.name == 'Symbol' {
		dump('type_sym')
		println(type_sym)
		println(type_sym.has_method(encode_json_member_name))
		println(type_sym.has_method('str'))
	}
	mut has_ser_json_method := false
	mut has_str_method := false
	for {
		if type_sym.has_method(encode_json_member_name) {
			has_ser_json_method = true
			break
		}
		if type_sym.has_method('str') {
			has_str_method = true
			break
		}
		info := type_sym.info
		if info is ast.Alias {
			type_sym = self.table.get_type_symbol(info.parent_type)
			$if debug {
				println(term.red(type_sym.name))
				dump(type_sym.name)
			}
		} else {
			break
		}
	}
	right := if typ == ast.string_type {
		field
	} else if has_ser_json_method {
		ast.Expr(ast.CallExpr{
			name: encode_json_member_name
			left: field
			scope: self.scope()
			is_method: true
		})
	} else if has_str_method {
		// print(field_name)
		_ = $if debug {
			dump(type_sym.name)
			true
		} $else {
			true
		}

		ast.Expr(ast.CallExpr{
			name: 'str'
			left: field
			scope: self.scope()
			is_method: true
		})
	} else {
		info := &type_sym.info
		match info {
			ast.Map {
				field
			}
			ast.Array {
				// $if debug {
				// 	dump(info)
				// }

				// elem_type_sym := self.table.get_type_symbol(type_sym.info.elem_type)
				
				// match elem_type_sym.info {

				// }
				j2any := self.find_type_or_add_placeholder('json2.Any', .v)
				ast.Expr(ast.CastExpr{
					typ: j2any
					expr: ast.CallExpr{
						name: 'map'
						args: [ast.CallArg {
							is_mut: false
							share: .mut_t
							expr: ast.CastExpr{
								typ: j2any
								expr: get_type_recursively(mut self, self.ident('it'), info.elem_type)
							}
						}]
						left: field
						scope: self.scope()
						is_method: true
					}
				})
			}
			ast.Enum {
				ast.Expr(ast.CallExpr{
					name: 'str'
					left: field
					scope: self.scope()
					is_method: true
				})
			}
			ast.Struct {
				ast.Expr(ast.CallExpr{
					name: encode_json_member_name
					left: field
					scope: self.scope()
					is_method: true
				})
			}
			else {
				field
			}
		}
	}
	return right
}


fn get_js_field_name(field ast.StructField) string {
	mut name := field.name
	for attr in field.attrs {
		if attr.name == 'json' {
			name = attr.arg
		}
		$if debug_attr ? {
			println(attr)
		}
	}
	return name
}
