module deser_json

import v.ast
import tool.codegen.util {str_to_type}
import tool.codegen.codegen {Codegen}

// generates
// ```vlang
// fn macro_decode_json__my_struct_name(j json2.Any) ?MyStructName { ... }
// ```
pub fn add_decode_json_fn(mut self Codegen, stmt ast.StructDecl) {
	// mut body_stmts := []ast.Stmt{}
	mut body_stmts := get_decode_json_base_stmts(mut self)

	body_stmts << ast.Return{
		exprs: [ast.Expr(ast.StructInit {
			// typ: self.table.get_type_symbol(self.table.type_idxs[stmt.name])
			typ: self.find_type_or_add_placeholder(stmt.name, .v)
			fields: stmt.fields.map(gen_struct_init_field(mut self, it))
			// fields: [
			// 	ast.StructInitField{
			// 		name: 'field_name'
			// 		expr: self.string_literal('a')
			// 	}
			// ]
		})]
	}
	mut params := [ast.Param{ name: 'j', typ: self.find_type_or_add_placeholder('json2.Any', .v) }]
	self.add_fn(name: get_decode_fn_name(stmt.name), return_type: ast.ovoid_type, body_stmts: body_stmts, params: params, comments: [
		self.gen_comment(text: 'generated by macro "derive_Deser')
		self.gen_comment(text: 'Example: ${decode_json_fn_name}<${stmt.name.split('.').last()}>(text)')
	])
}

fn get_struct_name_without_module(struct_name string) string {
	mut name := struct_name
	parts := name.split('.')

	if parts.len > 1 {
		name = parts[1]
	}
	return name
}
fn get_decode_fn_name(struct_name string) string {
	return '${decode_json_fn_name}__${to_snake_case(get_struct_name_without_module(struct_name))}'
}

fn get_decode_map_fn_name(struct_name string, depth int) string {
	mut res := '${decode_json_fn_name}__'
	for _ in 0..depth {
		res += 'map_'
	}
	name := get_struct_name_without_module(struct_name)
	res += '_${to_snake_case(name)}'
	return res
}
fn gen_struct_init_field(mut self Codegen, field ast.StructField) ast.StructInitField {
	return ast.StructInitField{
		name: field.name
		expr: get_assign_right_expr__fn(mut self, field.name, get_js_field_name(field), field.typ)
	}
}

fn get_map_depth(type_name string) int {
	mut temp := type_name
	mut depth := 0
	if temp.starts_with('map[string]') {
		
	}
}

fn get_assign_right_expr__fn(mut self Codegen, field_name string, js_field_name string, typ ast.Type) ast.Expr {
	if typ > ast.builtin_type_names.len {
		type_sym := self.table.get_type_symbol(typ)
		if type_sym.name.starts_with('map[string]') {
			// map
			// type_arg := type_sym.name.split_nth(']', 2)[1]

			type_arg := type_sym.name[10..]
			type_arg_idx := ast.Type(self.table.type_idxs[type_arg])
			return ast.Expr(ast.CallExpr{
					name: decode_json_map_fn_name
					args: [ast.CallArg {
						expr: ast.CallExpr{
							name: 'as_map'
							left: ast.IndexExpr{
								index: self.string_literal(js_field_name)
								left: self.ident(json2_map_name)
								or_expr: ast.OrExpr{ kind: .block, stmts: [self.integer_literal_stmt(0)] } // ast.CastExpr('json2.Any')
							}
							scope: self.scope(), is_method: true
						}
					}]
					concrete_types: [type_arg_idx]
					scope: self.scope(), is_method: false // left: self.ident('j')
					or_block: ast.OrExpr{ kind: .propagate }
			})
		} else if type_sym.name.starts_with('[') {
			// array
			type_arg := type_sym.name.split_nth(']', 2)[1]
			type_arg_idx := ast.Type(self.table.type_idxs[type_arg])
			return ast.Expr(ast.CallExpr{
					name: decode_json_array_fn_name
					args: [ast.CallArg {
						expr: ast.CallExpr{
							name: 'arr'
							left: ast.IndexExpr{
								index: self.string_literal(js_field_name)
								left: self.ident(json2_map_name)
								or_expr: ast.OrExpr{ kind: .block, stmts: [self.integer_literal_stmt(0)] }
							}
							scope: self.scope(), is_method: true
						}
					}]
					concrete_types: [type_arg_idx]
					scope: self.scope(), is_method: false // left: self.ident('j')
					or_block: ast.OrExpr{ kind: .propagate }
			})
		}
		// else {
			// 'json'
			mut decode_fn_name := decode_json_fn_name
			mut concrete_types := [typ]
			type_info := type_sym.info
			if type_info is ast.Enum {
				for attr in self.table.enum_decls[type_sym.name].attrs {
					if attr.name == 'deser_json_with' {
						decode_fn_name = attr.arg
						concrete_types.pop()
					}
				}
			}
			if type_info is ast.Struct {
				for attr in type_info.attrs {
					if attr.name == 'deser_json_with' {
						decode_fn_name = attr.arg
						concrete_types.pop()
					}
				}
			}
			return ast.Expr(ast.CallExpr{
					name: decode_fn_name
					args: [ast.CallArg {
						expr: ast.IndexExpr{
							index: self.string_literal(js_field_name)
							left: self.ident(json2_map_name)
							or_expr: ast.OrExpr{ kind: .block, stmts: [self.integer_literal_stmt(0)] }
						}
					}]
					concrete_types: concrete_types
					scope: self.scope(), is_method: false // left: self.ident('j')
					or_block: ast.OrExpr{ kind: .propagate }
				})
		// }
	} else if typ == ast.array_type_idx {
		return ast.Expr(ast.EmptyExpr{}) // TODO:
	} else if typ == ast.map_type_idx {
		return ast.Expr(ast.EmptyExpr{}) // TODO:
	} else {
		method_name, cast_type := get_json2_method_name(typ)
		mut expr := ast.Expr(ast.CallExpr{
				name: method_name
				left: ast.IndexExpr{
					index: self.string_literal(js_field_name)
					left: self.ident(json2_map_name)
					or_expr: ast.OrExpr{ kind: .block, stmts: [self.integer_literal_stmt(0)] }
				}
				scope: self.scope()
				is_method: true
			})
		if cast_type > 0 {
			return ast.CastExpr{
				typ: cast_type
				expr: expr
			}
		}
		return expr
	}
}
