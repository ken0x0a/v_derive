module ser

import v.ast { EnumDecl, Stmt, StructDecl, SumTypeDecl }
import v.token
import codegen { Codegen }
import common
import util { get_type_name_without_module }

// ```v
// pub fn (self Product) bin_encode(mut buf []byte) int {
// 	mut pos := 0
// 	pos += bincode.encode(mut buf, self.name)
// 	pos += bincode.encode(mut buf[pos..], self.desc)
// 	pos += bincode.encode(mut buf[pos..], self.inventory)
// 	pos += bincode.encode(mut buf[pos..], self.price)
// 	return pos
// }
// ```
pub fn add_encode_fn_for_struct(mut cg Codegen, decl StructDecl) {
	fn_name := common.fn_method_name_encode
	mut params := get_params(mut cg)
	return_type := ast.int_type

	mut body_stmts := []Stmt{cap: decl.fields.len + 2}
	body_stmts << base_assign_stmt(mut cg)
	for idx, field in decl.fields {
		body_stmts << gen_encode_and_plus_assign(mut cg, field, idx)
	}
	body_stmts << Stmt(ast.Return{
		exprs: [cg.ident(ident_name_encode_pos)]
	})
	cg.add_struct_method(
		struct_name: decl.name.split('.').last()
		is_mut: false
		name: fn_name
		return_type: return_type
		body_stmts: body_stmts
		params: params
		comments: [
			cg.gen_comment(text: 'generated by macro "$macro_name"'),
		]
	)
}

// ```v
// len += bincode.encode(mut b, self.a)
// ```
fn gen_encode_and_plus_assign(mut cg Codegen, field ast.StructField, idx int) ast.Stmt {
	field_sel := ast.SelectorExpr{ // 'self.$field'
		field_name: field.name
		expr: cg.ident(common.ident_name_self)
		scope: cg.scope()
	}

	arg1 := if idx == 0 {
		cg.ident(ident_name_bytes)
	} else {
		ast.Expr(ast.IndexExpr{
			left: cg.ident(ident_name_bytes)
			index: ast.RangeExpr{has_low: true, low: cg.ident(ident_name_encode_pos)}
		})
	}
	right := ast.Expr(ast.CallExpr{
		name: 'encode'
		left: cg.ident(common.mod_name)
		scope: cg.scope()
		is_method: true
		args: [
			ast.CallArg {expr: arg1, is_mut: true},
			ast.CallArg {expr: field_sel},
		]
	})
	return ast.AssignStmt{
		left: [cg.ident(ident_name_encode_pos)]
		right: [right]
		op: token.Kind.plus_assign
	}
}
